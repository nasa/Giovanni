netcdf ss.scrubbed.AIRX3STD_006_Temperature_A.20090119 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	TempPrsLvls_A = 24 ;
	lat = 2 ;
	lon = 2 ;
variables:
	float AIRX3STD_006_Temperature_A(time, TempPrsLvls_A, lat, lon) ;
		AIRX3STD_006_Temperature_A:_FillValue = -9999.f ;
		AIRX3STD_006_Temperature_A:standard_name = "air_temperature" ;
		AIRX3STD_006_Temperature_A:long_name = "Atmospheric Temperature Profile, 1000 to 1 hPa, daytime (ascending), AIRS, 1 x 1 deg." ;
		AIRX3STD_006_Temperature_A:units = "K" ;
		AIRX3STD_006_Temperature_A:missing_value = -9999.f ;
		AIRX3STD_006_Temperature_A:coordinates = "time TempPrsLvls_A lat lon" ;
		AIRX3STD_006_Temperature_A:quantity_type = "Air Temperature" ;
		AIRX3STD_006_Temperature_A:product_short_name = "AIRX3STD" ;
		AIRX3STD_006_Temperature_A:product_version = "006" ;
		AIRX3STD_006_Temperature_A:Serializable = "True" ;
	float TempPrsLvls_A(TempPrsLvls_A) ;
		TempPrsLvls_A:standard_name = "Pressure" ;
		TempPrsLvls_A:long_name = "Pressure Levels Temperature Profile, daytime (ascending) node" ;
		TempPrsLvls_A:units = "hPa" ;
		TempPrsLvls_A:positive = "down" ;
		TempPrsLvls_A:_CoordinateAxisType = "GeoZ" ;
	int dataday(time) ;
		dataday:standard_name = "Standardized Date Label" ;
	float lat(lat) ;
		lat:_FillValue = -9999.f ;
		lat:long_name = "Latitude" ;
		lat:missing_value = -9999.f ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
	float lon(lon) ;
		lon:_FillValue = -9999.f ;
		lon:long_name = "Longitude" ;
		lon:missing_value = -9999.f ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
	int time(time) ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00" ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:start_time = "2009-01-19T00:00:00Z" ;
		:end_time = "2009-01-19T23:59:59Z" ;
		:temporal_resolution = "daily" ;
		:nco_openmp_thread_number = 1 ;
		:NCO = "4.2.1" ;
		:history = "Mon Jul  1 13:59:57 2013: ncks -d lat,47.,49. -d lon,-148.,-146. scrubbed.AIRX3STD_006_Temperature_A.20090119.nc ss.scrubbed.AIRX3STD_006_Temperature_A.20090119.nc" ;
data:

 AIRX3STD_006_Temperature_A =
  277.25, 277.4375,
  277.5625, 276.5625,
  272.25, 272.75,
  272.5625, 271.4375,
  269.625, 270.4375,
  269.6875, 269.4375,
  262.9375, 263.1875,
  262.4375, 263.0625,
  253.8438, 253.9688,
  253.6875, 254.4062,
  244.1875, 244.1875,
  243.375, 243.625,
  234.5625, 234.3438,
  233.75, 233.5625,
  230.6562, 231.0625,
  231.0938, 231.2812,
  229.5, 230.5938,
  229.8438, 230.875,
  229.3438, 230.375,
  229.5312, 230.4062,
  226.0312, 226.25,
  226.2188, 226.4375,
  218.6875, 218.0625,
  219.375, 218.7188,
  217.125, 216.5625,
  217.7812, 216.8125,
  217.4688, 216.9375,
  217.5625, 216.7812,
  217.1562, 216.5312,
  216.9062, 216.5625,
  217.75, 217.0312,
  218.0312, 217.25,
  219.125, 218.375,
  219.6875, 218.5938,
  222.8125, 222.3125,
  223.5, 222.625,
  229.0938, 228.25,
  229.9688, 228.5,
  236.5938, 235.5,
  236.9688, 235.25,
  241.375, 240.625,
  240.0938, 239.7812,
  241.0312, 240.6562,
  239.0625, 239.5938,
  240.6875, 240.625,
  238.8125, 239.5,
  240.9688, 241.1562,
  239.8438, 240.4062 ;

 TempPrsLvls_A = 1000, 925, 850, 700, 600, 500, 400, 300, 250, 200, 150, 100, 
    70, 50, 30, 20, 15, 10, 7, 5, 3, 2, 1.5, 1 ;

 dataday = 2009019 ;

 lat = 47.5, 48.5 ;

 lon = -147.5, -146.5 ;

 time = 1232323200 ;
}
