netcdf t_nccorrelate_3d {
dimensions:
	longitude = 2 ;
	latitude = 2 ;
variables:
	double longitude(longitude) ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
		longitude:units = "degrees_east" ;
	double latitude(latitude) ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
		latitude:units = "degrees_north" ;
	double correlation(latitude, longitude) ;
		correlation:long_name = "correlation" ;
		correlation:_FillValue = 9.96920996838687e+36 ;
		correlation:quantity_type = "correlation" ;
	double slope(latitude, longitude) ;
		slope:long_name = "slope" ;
		slope:_FillValue = 9.96920996838687e+36 ;
	double offset(latitude, longitude) ;
		offset:long_name = "offset" ;
		offset:_FillValue = 9.96920996838687e+36 ;
	double time_matched_difference(latitude, longitude) ;
		time_matched_difference:long_name = "time_matched_difference" ;
		time_matched_difference:_FillValue = 9.96920996838687e+36 ;
		time_matched_difference:quantity_type = "difference" ;
	double sum_x(latitude, longitude) ;
		sum_x:long_name = "sum_x" ;
		sum_x:_FillValue = 9.96920996838687e+36 ;
	double sum_y(latitude, longitude) ;
		sum_y:long_name = "sum_y" ;
		sum_y:_FillValue = 9.96920996838687e+36 ;
	double sum_xy(latitude, longitude) ;
		sum_xy:long_name = "sum_xy" ;
		sum_xy:_FillValue = 0. ;
	double sum_x2(latitude, longitude) ;
		sum_x2:long_name = "sum_x2" ;
		sum_x2:_FillValue = 0. ;
	double sum_y2(latitude, longitude) ;
		sum_y2:long_name = "sum_y2" ;
		sum_y2:_FillValue = 0. ;
	int n_samples(latitude, longitude) ;
		n_samples:long_name = "Number of samples" ;
		n_samples:quantity_type = "count" ;
		n_samples:units = "count" ;

// global attributes:
		:Conventions = "CF-1.4" ;
data:

 longitude = -147.5, -146.5 ;

 latitude = 47.5, 48.5 ;

 correlation =
  0.983477394684323, 0.997048138338237,
  0.983479615753215, 0.995132631132934 ;

 slope =
  _, 0.939623558520744,
  _, 0.714959631698477 ;

 offset =
  43.6183148842875, 16.1008731719171,
  107.537036319516, 71.4619422533852 ;

 time_matched_difference =
  0.0520985921223958, -1.125,
  -0.0728708902994792, -0.635340372721354 ;

 sum_x =
  741.6875, 744.125,
  742.312591552734, 745.437591552734 ;

 sum_y =
  741.531204223633, 747.5,
  742.531204223633, 747.343612670898 ;

 sum_xy =
  183363.897870062, 185466.52734375,
  183768.292900085, 185752.768156047 ;

 sum_x2 =
  183410.209688191, 184632.9453125,
  183743.532007222, 185300.461957936 ;

 sum_y2 =
  183319.946698191, 186304.4296875,
  183806.541077616, 186212.73138333 ;

 n_samples =
  3, 3,
  3, 3 ;
}
