netcdf ss.scrubbed.AIRX3STD_006_Temperature_D.20090119 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	TempPrsLvls_D = 24 ;
	lat = 2 ;
	lon = 2 ;
variables:
	float AIRX3STD_006_Temperature_D(time, TempPrsLvls_D, lat, lon) ;
		AIRX3STD_006_Temperature_D:_FillValue = -9999.f ;
		AIRX3STD_006_Temperature_D:standard_name = "air_temperature" ;
		AIRX3STD_006_Temperature_D:long_name = "Atmospheric Temperature Profile, 1000 to 1 hPa, nighttime (descending), AIRS, 1 x 1 deg." ;
		AIRX3STD_006_Temperature_D:units = "K" ;
		AIRX3STD_006_Temperature_D:missing_value = -9999.f ;
		AIRX3STD_006_Temperature_D:coordinates = "time TempPrsLvls_D lat lon" ;
		AIRX3STD_006_Temperature_D:quantity_type = "Air Temperature" ;
		AIRX3STD_006_Temperature_D:product_short_name = "AIRX3STD" ;
		AIRX3STD_006_Temperature_D:product_version = "006" ;
		AIRX3STD_006_Temperature_D:Serializable = "True" ;
	float TempPrsLvls_D(TempPrsLvls_D) ;
		TempPrsLvls_D:standard_name = "Pressure" ;
		TempPrsLvls_D:long_name = "Pressure Levels Temperature Profile, nighttime (descending) node" ;
		TempPrsLvls_D:units = "hPa" ;
		TempPrsLvls_D:positive = "down" ;
		TempPrsLvls_D:_CoordinateAxisType = "GeoZ" ;
	int dataday(time) ;
		dataday:standard_name = "Standardized Date Label" ;
	float lat(lat) ;
		lat:_FillValue = -9999.f ;
		lat:long_name = "Latitude" ;
		lat:missing_value = -9999.f ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
	float lon(lon) ;
		lon:_FillValue = -9999.f ;
		lon:long_name = "Longitude" ;
		lon:missing_value = -9999.f ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
	int time(time) ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00" ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:start_time = "2009-01-19T00:00:00Z" ;
		:end_time = "2009-01-19T23:59:59Z" ;
		:temporal_resolution = "daily" ;
		:nco_openmp_thread_number = 1 ;
		:NCO = "4.2.1" ;
		:history = "Mon Jul  1 13:59:57 2013: ncks -d lat,47.,49. -d lon,-148.,-146. scrubbed.AIRX3STD_006_Temperature_D.20090119.nc ss.scrubbed.AIRX3STD_006_Temperature_D.20090119.nc" ;
data:

 AIRX3STD_006_Temperature_D =
  277.1875, 277.9375,
  277.5625, 277.125,
  271.875, 272.5625,
  272.375, 272.0625,
  269.625, 269.9375,
  270.3125, 269.8125,
  262.6875, 263.0625,
  263.25, 263.1875,
  254.125, 254.9688,
  254.4688, 254.9688,
  244, 245.1875,
  244.6562, 245.2812,
  233.375, 234.5,
  234.1562, 235,
  231.2188, 231.9375,
  231.2188, 232.0312,
  232.1562, 232.9688,
  231.7812, 232.4688,
  231.8438, 232.2812,
  231.4688, 231.7188,
  227.2188, 226.625,
  226.9062, 226.4375,
  219.25, 218.25,
  219.3125, 218.4375,
  217.9062, 217.3438,
  218.4688, 217.75,
  217.9062, 217.375,
  218.0938, 217.6875,
  218.2812, 217.5625,
  218.2188, 217.6562,
  218.4062, 218.0625,
  218.1875, 217.75,
  218.875, 218.7812,
  218.8438, 218.375,
  223.2188, 223.2188,
  223.0938, 222.5,
  230.0625, 230.0625,
  229.6875, 229.125,
  239.1875, 238.8125,
  238.5312, 237.9375,
  247.8125, 245.6875,
  247.1562, 246,
  247.4688, 245.375,
  247.125, 246.25,
  245.0625, 243.2812,
  244.8125, 244.0625,
  240.875, 239.9688,
  240.6875, 240.2812 ;

 TempPrsLvls_D = 1000, 925, 850, 700, 600, 500, 400, 300, 250, 200, 150, 100, 
    70, 50, 30, 20, 15, 10, 7, 5, 3, 2, 1.5, 1 ;

 dataday = 2009019 ;

 lat = 47.5, 48.5 ;

 lon = -147.5, -146.5 ;

 time = 1232323200 ;
}
