netcdf AIRS_Temp_D.20090118.500hPa {
dimensions:
	time = UNLIMITED ; // (1 currently)
	TempPrsLvls_D = 1 ;
	lat = 2 ;
	lon = 2 ;
variables:
	float AIRX3STD_006_Temperature_D(time, TempPrsLvls_D, lat, lon) ;
		AIRX3STD_006_Temperature_D:_FillValue = -9999.f ;
		AIRX3STD_006_Temperature_D:standard_name = "air_temperature" ;
		AIRX3STD_006_Temperature_D:long_name = "Atmospheric Temperature Profile, 1000 to 1 hPa, nighttime (descending), AIRS, 1 x 1 deg." ;
		AIRX3STD_006_Temperature_D:units = "K" ;
		AIRX3STD_006_Temperature_D:missing_value = -9999.f ;
		AIRX3STD_006_Temperature_D:coordinates = "time TempPrsLvls_D lat lon" ;
		AIRX3STD_006_Temperature_D:quantity_type = "Air Temperature" ;
		AIRX3STD_006_Temperature_D:product_short_name = "AIRX3STD" ;
		AIRX3STD_006_Temperature_D:product_version = "006" ;
		AIRX3STD_006_Temperature_D:Serializable = "True" ;
	float TempPrsLvls_D(TempPrsLvls_D) ;
		TempPrsLvls_D:standard_name = "Pressure" ;
		TempPrsLvls_D:long_name = "Pressure Levels Temperature Profile, nighttime (descending) node" ;
		TempPrsLvls_D:units = "hPa" ;
		TempPrsLvls_D:positive = "down" ;
		TempPrsLvls_D:_CoordinateAxisType = "GeoZ" ;
	int dataday(time) ;
		dataday:standard_name = "Standardized Date Label" ;
	float lat(lat) ;
		lat:_FillValue = -9999.f ;
		lat:long_name = "Latitude" ;
		lat:missing_value = -9999.f ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
	float lon(lon) ;
		lon:_FillValue = -9999.f ;
		lon:long_name = "Longitude" ;
		lon:missing_value = -9999.f ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
	int time(time) ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00" ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:start_time = "2009-01-18T00:00:00Z" ;
		:end_time = "2009-01-18T23:59:59Z" ;
		:temporal_resolution = "daily" ;
		:nco_openmp_thread_number = 1 ;
		:NCO = "4.2.2" ;
		:history = "Thu Jul  4 19:19:54 2013: ncks -d TempPrsLvls_D,500.,500. AIRS_Temp_D.20090118.nc AIRS_Temp_D.20090118.500hPa.nc\n",
			"Mon Jul  1 13:59:57 2013: ncks -d lat,47.,49. -d lon,-148.,-146. scrubbed.AIRX3STD_006_Temperature_D.20090118.nc ss.scrubbed.AIRX3STD_006_Temperature_D.20090118.nc" ;
data:

 AIRX3STD_006_Temperature_D =
  246, 247.375,
  246.6875, 248.1562 ;

 TempPrsLvls_D = 500 ;

 dataday = 2009018 ;

 lat = 47.5, 48.5 ;

 lon = -147.5, -146.5 ;

 time = 1232236800 ;
}
