netcdf t_accumulate_1 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	Latitude = 8 ;
	Longitude = 3 ;
variables:
	int time(time) ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00" ;
	short Optical_Depth_Land_And_Ocean_Mean(time, Latitude, Longitude) ;
		Optical_Depth_Land_And_Ocean_Mean:coordinates = "time Latitude Longitude" ;
		Optical_Depth_Land_And_Ocean_Mean:Level_2_Pixel_Values_Read_As = "Real" ;
		Optical_Depth_Land_And_Ocean_Mean:Quality_Assurance_Data_Set = "None" ;
		Optical_Depth_Land_And_Ocean_Mean:Derived_From_Level_2_Data_Set = "Optical_Depth_Land_And_Ocean" ;
		Optical_Depth_Land_And_Ocean_Mean:long_name = "Aerosol Optical Thickness at 0.55 microns for both Ocean (best) and Land (corrected): Mean" ;
		Optical_Depth_Land_And_Ocean_Mean:valid_range = -100s, 5000s ;
		Optical_Depth_Land_And_Ocean_Mean:Included_Level_2_Nighttime_Data = "False" ;
		Optical_Depth_Land_And_Ocean_Mean:Aggregation_Data_Set = "None" ;
		Optical_Depth_Land_And_Ocean_Mean:_FillValue = -9999s ;
		Optical_Depth_Land_And_Ocean_Mean:Statistic_Type = "Simple" ;
		Optical_Depth_Land_And_Ocean_Mean:add_offset = 0. ;
		Optical_Depth_Land_And_Ocean_Mean:units = "1" ;
		Optical_Depth_Land_And_Ocean_Mean:scale_factor = 0.001 ;
		Optical_Depth_Land_And_Ocean_Mean:quantity_type = "Aerosol Optical Depth" ;
	double Latitude(Latitude) ;
		Latitude:long_name = "Latitude" ;
		Latitude:units = "degrees_north" ;
	double Longitude(Longitude) ;
		Longitude:long_name = "Longitude" ;
		Longitude:units = "degrees_east" ;

// global attributes:
		:Conventions = "CF-1.4" ;
data:

 time = 1262217600 ;

 Optical_Depth_Land_And_Ocean_Mean =
  _, _, 314,
  475, 300, 420,
  515, 498, 482,
  564, 502, 415,
  650, 492, 434,
  676, 626, _,
  707, 632, 337,
  _, 329, 377 ;

 Latitude = 34.5, 33.5, 32.5, 31.5, 30.5, 29.5, 28.5, 27.5 ;

 Longitude = 116.5, 117.5, 118.5 ;
}
